Bit#(32) compileTime = 1278088049; // Verilog Fri Jul 2 12:27:29 EDT 2010
