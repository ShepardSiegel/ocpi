Bit#(32) compileTime = 1314223867; // Verilog Wed Aug 24 18:11:07 EDT 2011
