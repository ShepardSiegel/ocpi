Bit#(32) compileTime = 1275592252; // Verilog Thu Jun 3 15:10:52 EDT 2010
