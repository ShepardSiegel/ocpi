Bit#(32) compileTime = 1277891087; // Verilog Wed Jun 30 05:44:47 EDT 2010
