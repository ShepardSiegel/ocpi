// OCTG.bsv
// Copyright (c) 2009 Atomic Rules LLC - ALL RIGHTS RESERVED

package OCTG;

import OCTG_nosm::*;
import OCTG_genchk::*;
import OCTG_dmaFP::*;
import OCTG_dmaFC::*;
import OCTG_dma2push::*;

export OCTG_nosm::*;
export OCTG_genchk::*;
export OCTG_dmaFP::*;
export OCTG_dmaFC::*;
export OCTG_dma2push::*;

endpackage: OCTG
