Bit#(32) compileTime = 1276725574; // Verilog Wed Jun 16 17:59:34 EDT 2010
