Bit#(32) compileTime = 1304974432; // Verilog Mon May 9 16:53:52 EDT 2011
