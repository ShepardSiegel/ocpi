Bit#(32) compileTime = 1317476396; // Verilog Sat Oct 1 09:39:56 EDT 2011
