Bit#(32) compileTime = 1289939306; // Verilog Tue Nov 16 15:28:26 EST 2010
