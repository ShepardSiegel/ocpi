Bit#(32) compileTime = 1275387336; // Verilog Tue Jun 1 06:15:36 EDT 2010
