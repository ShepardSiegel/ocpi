Bit#(32) compileTime = 1277736309; // ISim Mon Jun 28 10:45:09 EDT 2010
