Bit#(32) compileTime = 1289150389; // Verilog Sun Nov 7 12:19:49 EST 2010
