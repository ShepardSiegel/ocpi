Bit#(32) compileTime = 1284043682; // Verilog Thu Sep 9 10:48:02 EDT 2010
