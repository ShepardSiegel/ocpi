Bit#(32) compileTime = 1285680713; // Verilog Tue Sep 28 09:31:53 EDT 2010
