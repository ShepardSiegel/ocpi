Bit#(32) compileTime = 1277994263; // Verilog Thu Jul 1 10:24:23 EDT 2010
