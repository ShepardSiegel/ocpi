Bit#(32) compileTime = 1293105349; // Verilog Thu Dec 23 06:55:49 EST 2010
