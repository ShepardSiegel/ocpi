Bit#(32) compileTime = 1383602750; // Verilog Mon Nov 4 17:05:50 EST 2013
