Bit#(32) compileTime = 1295883839; // Verilog Mon Jan 24 10:43:59 EST 2011
