Bit#(32) compileTime = 1278606896; // Verilog Thu Jul 8 12:34:56 EDT 2010
