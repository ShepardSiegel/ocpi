// DelayAssy.bsv
// Copyright (c) 2010 Atomic Rules LLC - ALL RIGHTS RESERVED
//
// This is a human-generated BSV source file based upon the provided "delayAssy_defs.v"
// It is intended to be a guide and template towards OpenCPI's programatic generation of this file
// this may be called "OpenCPI exportCPI for BSV"


package DelayAssy; // Name this package 

import OCWip::*;     // Include the OpenCPI BSV WIP package 
import Vector::*;    // Include the Bluespec Vector package

// Local typedefs that specialize the various interaces to a shorthand
// Theses type paramaters are derrived from WIP attributes
// Autogenerated comments should include workername that use these types
// We use the I_ prefix for interface Types so that names have no case restrictions
typedef WciEs                    I_wci0;    // describe WIP attributes here
typedef WciEs                    I_wci1;    // describe WIP attributes here
typedef WciEs                    I_wci2;    // describe WIP attributes here
typedef Wmemi_Em#(36,12,128,16)  I_wmemi0;  // describe WIP attributes here
typedef Wsi_Es#(12,32,4,8,1)     I_adc;     // describe WIP attributes here
typedef Wsi_Em#(12,32,4,8,1)     I_dac;     // describe WIP attributes here
typedef Wmi_Em#(14,12,32,0,0,32) I_FC;      // describe WIP attributes here
typedef Wmi_Em#(14,12,32,0,0,32) I_FP;      // describe WIP attributes here

// Define the interface for a thin Verilog wrapper around the assemply code
// Name the interface as the concatenation of V, package_name, Ifc
// We use the i_ prefix for sub-interface instance names so that names have no case restrictions
// Autogenerated comments should include real workernames...
interface VDelayAssyIfc;
  interface I_wci0   i_wci0;      // WCI Slave  Interface 0 for worker workername
  interface I_wci1   i_wci1;      // WCI Slave  Interface 1 for worker workername
  interface I_wci2   i_wci2;      // WCI Slave  Interface 2 for worker workername
  interface I_wmemi0 i_wmemi0;    // WMemi Master Interface supporting worker workername
  interface I_adc    i_adc;       // WSI Slave  interfcae from ADC to worker workername
  interface I_dac    i_dac;       // WSI Master interfcae from worker workername to DAC
  interface I_FC     i_FC;        // WMI Master interface for worker workername
  interface I_FP     i_FP;        // WMI Master interface for worker workername
endinterface: VDelayAssyIfc

// Use importBVI to bind the signal names in the underlying Verilog to BSV methods
import "BVI" delayAssy_defs =
module vMkDelayAssy#(Clock wciClk, Vector#(3,Reset) wciRst) (VDelayAssyIfc);

  default_clock no_clock;
  default_reset no_reset;
  input_clock   wciClk (wci_Clk)   = wciClk;  // The common clock used for all WCI Slaves in the assembly
  input_reset   wciRst0(wci0_MReset_n)  = wciRst[0];
  input_reset   wciRst1(wci1_MReset_n)  = wciRst[1];
  input_reset   wciRst2(wci2_MReset_n)  = wciRst[2];

// For each sub-interface, list all the Action and Value methods and their unique associated Verilog signals...

interface I_wci0 i_wci0;
  method mCmd       (wci0_MCmd)        enable((*inhigh*)en0)   clocked_by(wciClk) reset_by(wciRst0);        
  method mAddrSpace (wci0_MAddrSpace)  enable((*inhigh*)en1)   clocked_by(wciClk) reset_by(wciRst0);        
  method mByteEn    (wci0_MByteEn)     enable((*inhigh*)en2)   clocked_by(wciClk) reset_by(wciRst0);        
  method mAddr      (wci0_MAddr)       enable((*inhigh*)en3)   clocked_by(wciClk) reset_by(wciRst0);        
  method mData      (wci0_MData)       enable((*inhigh*)en4)   clocked_by(wciClk) reset_by(wciRst0);        
  method mFlag      (wci0_MFlag)       enable((*inhigh*)en5)   clocked_by(wciClk) reset_by(wciRst0);        
  method wci0_SResp       sResp                                clocked_by(wciClk) reset_by(wciRst0);        
  method wci0_SData       sData                                clocked_by(wciClk) reset_by(wciRst0);        
  method wci0_SThreadBusy sThreadBusy                          clocked_by(wciClk) reset_by(wciRst0);        
  method wci0_SFlag       sFlag                                clocked_by(wciClk) reset_by(wciRst0);        
endinterface: i_wci0

interface I_wci1 i_wci1;
  method mCmd       (wci1_MCmd)        enable((*inhigh*)en6)   clocked_by(wciClk) reset_by(wciRst1);        
  method mAddrSpace (wci1_MAddrSpace)  enable((*inhigh*)en7)   clocked_by(wciClk) reset_by(wciRst1);        
  method mByteEn    (wci1_MByteEn)     enable((*inhigh*)en8)   clocked_by(wciClk) reset_by(wciRst1);        
  method mAddr      (wci1_MAddr)       enable((*inhigh*)en9)   clocked_by(wciClk) reset_by(wciRst1);        
  method mData      (wci1_MData)       enable((*inhigh*)en10)  clocked_by(wciClk) reset_by(wciRst1);        
  method mFlag      (wci1_MFlag)       enable((*inhigh*)en11)  clocked_by(wciClk) reset_by(wciRst1);        
  method wci1_SResp       sResp                                clocked_by(wciClk) reset_by(wciRst1);        
  method wci1_SData       sData                                clocked_by(wciClk) reset_by(wciRst1);        
  method wci1_SThreadBusy sThreadBusy                          clocked_by(wciClk) reset_by(wciRst1);        
  method wci1_SFlag       sFlag                                clocked_by(wciClk) reset_by(wciRst1);        
endinterface: i_wci1

interface I_wci2 i_wci2;
  method mCmd       (wci2_MCmd)        enable((*inhigh*)en12)  clocked_by(wciClk) reset_by(wciRst2);        
  method mAddrSpace (wci2_MAddrSpace)  enable((*inhigh*)en13)  clocked_by(wciClk) reset_by(wciRst2);        
  method mByteEn    (wci2_MByteEn)     enable((*inhigh*)en14)  clocked_by(wciClk) reset_by(wciRst2);        
  method mAddr      (wci2_MAddr)       enable((*inhigh*)en15)  clocked_by(wciClk) reset_by(wciRst2);        
  method mData      (wci2_MData)       enable((*inhigh*)en16)  clocked_by(wciClk) reset_by(wciRst2);        
  method mFlag      (wci2_MFlag)       enable((*inhigh*)en17)  clocked_by(wciClk) reset_by(wciRst2);        
  method wci2_SResp       sResp                                clocked_by(wciClk) reset_by(wciRst2);        
  method wci2_SData       sData                                clocked_by(wciClk) reset_by(wciRst2);        
  method wci2_SThreadBusy sThreadBusy                          clocked_by(wciClk) reset_by(wciRst2);        
  method wci2_SFlag       sFlag                                clocked_by(wciClk) reset_by(wciRst2);        
endinterface: i_wci2

interface I_wmemi0 i_wmemi0;
  method sResp           (wmemi0_SResp)           enable((*inhigh*)en18) clocked_by(wciClk) reset_by(no_reset);
  method sRespLast       ()                     enable(wmemi0_SRespLast) clocked_by(wciClk) reset_by(no_reset);
  method sData           (wmemi0_SData)           enable((*inhigh*)en20) clocked_by(wciClk) reset_by(no_reset);
  method sCmdAccept      ()                    enable(wmemi0_SCmdAccept) clocked_by(wciClk) reset_by(no_reset);
  method sDataAccept     ()                   enable(wmemi0_SDataAccept) clocked_by(wciClk) reset_by(no_reset);
  method wmemi0_MCmd         mCmd                                        clocked_by(wciClk) reset_by(no_reset);
  method wmemi0_MReqLast     mReqLast                                    clocked_by(wciClk) reset_by(no_reset);
  method wmemi0_MAddr        mAddr                                       clocked_by(wciClk) reset_by(no_reset);
  method wmemi0_MBurstLength mBurstLength                                clocked_by(wciClk) reset_by(no_reset);
  method wmemi0_MDataValid   mDataValid                                  clocked_by(wciClk) reset_by(no_reset);
  method wmemi0_MDataLast    mDataLast                                   clocked_by(wciClk) reset_by(no_reset);
  method wmemi0_MData        mData                                       clocked_by(wciClk) reset_by(no_reset);
  method wmemi0_MDataByteEn  mDataByteEn                                 clocked_by(wciClk) reset_by(no_reset);
  method wmemi0_MReset_n     mReset_n                                    clocked_by(wciClk) reset_by(no_reset);
endinterface: i_wmemi0

interface I_adc i_adc;
  method mCmd          (adc_MCmd)           enable((*inhigh*)en25) clocked_by(wciClk) reset_by(no_reset);
  method mReqLast      ()                     enable(adc_MReqLast) clocked_by(wciClk) reset_by(no_reset);
  method mBurstPrecise ()                enable(adc_MBurstPrecise) clocked_by(wciClk) reset_by(no_reset);
  method mBurstLength  (adc_MBurstLength)   enable((*inhigh*)en28) clocked_by(wciClk) reset_by(no_reset);
  method mData         (adc_MData)          enable((*inhigh*)en29) clocked_by(wciClk) reset_by(no_reset);
  method mByteEn       (adc_MByteEn)        enable((*inhigh*)en30) clocked_by(wciClk) reset_by(no_reset);
  method mReqInfo      (adc_MReqInfo)       enable((*inhigh*)en31) clocked_by(wciClk) reset_by(no_reset);
  method mDataInfo     (adc_MDataInfo)      enable((*inhigh*)en32) clocked_by(wciClk) reset_by(no_reset);
  method mReset_n     ()                      enable(adc_MReset_n) clocked_by(wciClk) reset_by(no_reset);
  method adc_SThreadBusy sThreadBusy                               clocked_by(wciClk) reset_by(no_reset);
  method adc_SReset_n    sReset_n                                  clocked_by(wciClk) reset_by(no_reset);
endinterface: i_adc

interface I_dac i_dac;
  method sThreadBusy ()                    enable(dac_SThreadBusy) clocked_by(wciClk) reset_by(no_reset);
  method sReset_n    ()                       enable(dac_SReset_n) clocked_by(wciClk) reset_by(no_reset);
  method dac_MCmd          mCmd                                    clocked_by(wciClk) reset_by(no_reset);
  method dac_MReqLast      mReqLast                                clocked_by(wciClk) reset_by(no_reset);
  method dac_MBurstPrecise mBurstPrecise                           clocked_by(wciClk) reset_by(no_reset);
  method dac_MBurstLength  mBurstLength                            clocked_by(wciClk) reset_by(no_reset);
  method dac_MData         mData                                   clocked_by(wciClk) reset_by(no_reset);
  method dac_MByteEn       mByteEn                                 clocked_by(wciClk) reset_by(no_reset);
  method dac_MReqInfo      mReqInfo                                clocked_by(wciClk) reset_by(no_reset);
  method dac_MDataInfo     mDataInfo                               clocked_by(wciClk) reset_by(no_reset);
  method dac_MReset_n      mReset_n                                clocked_by(wciClk) reset_by(no_reset);
endinterface: i_dac

interface I_FC i_FC;
  method sResp           (FC_SResp)            enable((*inhigh*)en36) clocked_by(wciClk) reset_by(no_reset);
  method sData           (FC_SData)            enable((*inhigh*)en37) clocked_by(wciClk) reset_by(no_reset);
  method sThreadBusy     ()                    enable(FC_SThreadBusy) clocked_by(wciClk) reset_by(no_reset);
  method sDataThreadBusy ()                enable(FC_SDataThreadBusy) clocked_by(wciClk) reset_by(no_reset);
  method sFlag           (FC_SFlag)            enable((*inhigh*)en40) clocked_by(wciClk) reset_by(no_reset);
  method sReset_n        ()                       enable(FC_SReset_n) clocked_by(wciClk) reset_by(no_reset);
  method FC_MCmd         mCmd                                         clocked_by(wciClk) reset_by(no_reset);
  method FC_MReqLast     mReqLast                                     clocked_by(wciClk) reset_by(no_reset);
  method FC_MReqInfo     mReqInfo                                     clocked_by(wciClk) reset_by(no_reset);
  method FC_MAddrSpace   mAddrSpace                                   clocked_by(wciClk) reset_by(no_reset);
  method FC_MAddr        mAddr                                        clocked_by(wciClk) reset_by(no_reset);
  method FC_MBurstLength mBurstLength                                 clocked_by(wciClk) reset_by(no_reset);
  method FC_MDataValid   mDataValid                                   clocked_by(wciClk) reset_by(no_reset);
  method FC_MDataLast    mDataLast                                    clocked_by(wciClk) reset_by(no_reset);
  method FC_MData        mData                                        clocked_by(wciClk) reset_by(no_reset);
  method FC_MDataInfo    mDataInfo                                    clocked_by(wciClk) reset_by(no_reset);
  method FC_MDataByteEn  mDataByteEn                                  clocked_by(wciClk) reset_by(no_reset);
  method FC_MFlag        mFlag                                        clocked_by(wciClk) reset_by(no_reset);
  method FC_MReset_n     mReset_n                                     clocked_by(wciClk) reset_by(no_reset);
endinterface: i_FC

interface I_FP i_FP;
  method sResp           (FP_SResp)            enable((*inhigh*)en42) clocked_by(wciClk) reset_by(no_reset);
  method sData           (FP_SData)            enable((*inhigh*)en43) clocked_by(wciClk) reset_by(no_reset);
  method sThreadBusy     ()                    enable(FP_SThreadBusy) clocked_by(wciClk) reset_by(no_reset);
  method sDataThreadBusy ()                enable(FP_SDataThreadBusy) clocked_by(wciClk) reset_by(no_reset);
  method sFlag           (FP_SFlag)            enable((*inhigh*)en46) clocked_by(wciClk) reset_by(no_reset);
  method sReset_n        ()                       enable(FP_SReset_n) clocked_by(wciClk) reset_by(no_reset);
  method FP_MCmd         mCmd                                         clocked_by(wciClk) reset_by(no_reset);
  method FP_MReqLast     mReqLast                                     clocked_by(wciClk) reset_by(no_reset);
  method FP_MReqInfo     mReqInfo                                     clocked_by(wciClk) reset_by(no_reset);
  method FP_MAddrSpace   mAddrSpace                                   clocked_by(wciClk) reset_by(no_reset);
  method FP_MAddr        mAddr                                        clocked_by(wciClk) reset_by(no_reset);
  method FP_MBurstLength mBurstLength                                 clocked_by(wciClk) reset_by(no_reset);
  method FP_MDataValid   mDataValid                                   clocked_by(wciClk) reset_by(no_reset);
  method FP_MDataLast    mDataLast                                    clocked_by(wciClk) reset_by(no_reset);
  method FP_MData        mData                                        clocked_by(wciClk) reset_by(no_reset);
  method FP_MDataInfo    mDataInfo                                    clocked_by(wciClk) reset_by(no_reset);
  method FP_MDataByteEn  mDataByteEn                                  clocked_by(wciClk) reset_by(no_reset);
  method FP_MFlag        mFlag                                        clocked_by(wciClk) reset_by(no_reset);
  method FP_MReset_n     mReset_n                                     clocked_by(wciClk) reset_by(no_reset);
endinterface: i_FP

schedule
  ( i_wci0_mCmd, i_wci0_mAddrSpace, i_wci0_mByteEn, i_wci0_mAddr, i_wci0_mData, i_wci0_mFlag, i_wci0_sResp, i_wci0_sData, i_wci0_sThreadBusy, i_wci0_sFlag, i_wci1_mCmd, i_wci1_mAddrSpace, i_wci1_mByteEn, i_wci1_mAddr, i_wci1_mData, i_wci1_mFlag, i_wci1_sResp, i_wci1_sData, i_wci1_sThreadBusy, i_wci1_sFlag, i_wci2_mCmd, i_wci2_mAddrSpace, i_wci2_mByteEn, i_wci2_mAddr, i_wci2_mData, i_wci2_mFlag, i_wci2_sResp, i_wci2_sData, i_wci2_sThreadBusy, i_wci2_sFlag, 
  i_wmemi0_sResp, i_wmemi0_sRespLast, i_wmemi0_sData , i_wmemi0_sCmdAccept , i_wmemi0_sDataAccept , i_wmemi0_mCmd, i_wmemi0_mReqLast, i_wmemi0_mAddr, i_wmemi0_mBurstLength, i_wmemi0_mDataValid, i_wmemi0_mDataLast, i_wmemi0_mData, i_wmemi0_mDataByteEn, i_wmemi0_mReset_n,
  i_adc_mCmd , i_adc_mReqLast, i_adc_mBurstPrecise, i_adc_mBurstLength, i_adc_mData, i_adc_mByteEn, i_adc_mReqInfo , i_adc_mDataInfo, i_adc_mReset_n, i_adc_sThreadBusy, i_adc_sReset_n, i_dac_mCmd , i_dac_mReqLast, i_dac_mBurstPrecise, i_dac_mBurstLength, i_dac_mData, i_dac_mByteEn, i_dac_mReqInfo , i_dac_mDataInfo, i_dac_mReset_n, i_dac_sThreadBusy, i_dac_sReset_n, 
  i_FC_mCmd, i_FC_mReqLast, i_FC_mReqInfo, i_FC_mAddrSpace , i_FC_mAddr, i_FC_mBurstLength, i_FC_mDataValid, i_FC_mDataLast , i_FC_mData , i_FC_mDataInfo , i_FC_mDataByteEn, i_FC_mFlag, i_FC_mReset_n, i_FC_sResp, i_FC_sData, i_FC_sThreadBusy, i_FC_sDataThreadBusy, i_FC_sFlag , i_FC_sReset_n, i_FP_mCmd, i_FP_mReqLast, i_FP_mReqInfo, i_FP_mAddrSpace , i_FP_mAddr, i_FP_mBurstLength, i_FP_mDataValid, i_FP_mDataLast , i_FP_mData , i_FP_mDataInfo , i_FP_mDataByteEn, i_FP_mFlag, i_FP_mReset_n, i_FP_sResp, i_FP_sData, i_FP_sThreadBusy, i_FP_sDataThreadBusy, i_FP_sFlag , i_FP_sReset_n )
  CF
  ( i_wci0_mCmd, i_wci0_mAddrSpace, i_wci0_mByteEn, i_wci0_mAddr, i_wci0_mData, i_wci0_mFlag, i_wci0_sResp, i_wci0_sData, i_wci0_sThreadBusy, i_wci0_sFlag, i_wci1_mCmd, i_wci1_mAddrSpace, i_wci1_mByteEn, i_wci1_mAddr, i_wci1_mData, i_wci1_mFlag, i_wci1_sResp, i_wci1_sData, i_wci1_sThreadBusy, i_wci1_sFlag, i_wci2_mCmd, i_wci2_mAddrSpace, i_wci2_mByteEn, i_wci2_mAddr, i_wci2_mData, i_wci2_mFlag, i_wci2_sResp, i_wci2_sData, i_wci2_sThreadBusy, i_wci2_sFlag, 
  i_wmemi0_sResp, i_wmemi0_sRespLast, i_wmemi0_sData , i_wmemi0_sCmdAccept , i_wmemi0_sDataAccept , i_wmemi0_mCmd, i_wmemi0_mReqLast, i_wmemi0_mAddr, i_wmemi0_mBurstLength, i_wmemi0_mDataValid, i_wmemi0_mDataLast, i_wmemi0_mData, i_wmemi0_mDataByteEn, i_wmemi0_mReset_n,
  i_adc_mCmd , i_adc_mReqLast, i_adc_mBurstPrecise, i_adc_mBurstLength, i_adc_mData, i_adc_mByteEn, i_adc_mReqInfo , i_adc_mDataInfo, i_adc_mReset_n, i_adc_sThreadBusy, i_adc_sReset_n, i_dac_mCmd , i_dac_mReqLast, i_dac_mBurstPrecise, i_dac_mBurstLength, i_dac_mData, i_dac_mByteEn, i_dac_mReqInfo , i_dac_mDataInfo, i_dac_mReset_n, i_dac_sThreadBusy, i_dac_sReset_n, 
  i_FC_mCmd, i_FC_mReqLast, i_FC_mReqInfo, i_FC_mAddrSpace , i_FC_mAddr, i_FC_mBurstLength, i_FC_mDataValid, i_FC_mDataLast , i_FC_mData , i_FC_mDataInfo , i_FC_mDataByteEn, i_FC_mFlag, i_FC_mReset_n, i_FC_sResp, i_FC_sData, i_FC_sThreadBusy, i_FC_sDataThreadBusy, i_FC_sFlag , i_FC_sReset_n, i_FP_mCmd, i_FP_mReqLast, i_FP_mReqInfo, i_FP_mAddrSpace , i_FP_mAddr, i_FP_mBurstLength, i_FP_mDataValid, i_FP_mDataLast , i_FP_mData , i_FP_mDataInfo , i_FP_mDataByteEn, i_FP_mFlag, i_FP_mReset_n, i_FP_sResp, i_FP_sData, i_FP_sThreadBusy, i_FP_sDataThreadBusy, i_FP_sFlag , i_FP_sReset_n);

endmodule: vMkDelayAssy


// Make a synthesizable Verilog module out of our wrapper...
(* synthesize, no_default_clock, no_default_reset, clock_prefix="", reset_prefix="" *)
(* doc= "Place generated documenantion here. Ok to use\nto put data on the next line\nand the next" *)
module mkDelayAssy#(Clock wciClk, Vector#(3,Reset) wciRst) (VDelayAssyIfc);
  (* hide *)
  let _ifc <- vMkDelayAssy(wciClk, wciRst);
  return _ifc;
endmodule: mkDelayAssy

endpackage: DelayAssy

