Bit#(32) compileTime = 1283883897; // Verilog Tue Sep 7 14:24:57 EDT 2010
