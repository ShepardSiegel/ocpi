Bit#(32) compileTime = 1289854433; // Verilog Mon Nov 15 15:53:53 EST 2010
