Bit#(32) compileTime = 1277981370; // Verilog Thu Jul 1 06:49:30 EDT 2010
