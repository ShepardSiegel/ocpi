Bit#(32) compileTime = 1390764368; // Verilog Sun Jan 26 14:26:08 EST 2014
