Bit#(32) compileTime = 1277134387; // Verilog Mon Jun 21 11:33:07 EDT 2010
