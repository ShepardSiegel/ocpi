Bit#(32) compileTime = 1328629586; // Verilog Tue Feb 7 10:46:26 EST 2012
