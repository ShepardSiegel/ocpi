Bit#(32) compileTime = 1305398449; // Verilog Sat May 14 14:40:49 EDT 2011
