Bit#(32) compileTime = 1304970059; // Verilog Mon May 9 15:40:59 EDT 2011
