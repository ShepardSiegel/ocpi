Bit#(32) compileTime = 1308673301; // Verilog Tue Jun 21 12:21:41 EDT 2011
