Bit#(32) compileTime = 1281623583; // Verilog Thu Aug 12 10:33:03 EDT 2010
