Bit#(32) compileTime = 1297262873; // Bluesim Wed Feb 9 09:47:53 EST 2011
