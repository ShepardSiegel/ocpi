Bit#(32) compileTime = 1278970800; // Verilog Mon Jul 12 17:40:00 EDT 2010
