Bit#(32) compileTime = 1277336883; // Verilog Wed Jun 23 19:48:03 EDT 2010
