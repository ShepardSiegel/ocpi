Bit#(32) compileTime = 1289236835; // Verilog Mon Nov 8 12:20:35 EST 2010
