Bit#(32) compileTime = 1282567602; // Verilog Mon Aug 23 08:46:42 EDT 2010
