Bit#(32) compileTime = 1314315997; // Verilog Thu Aug 25 19:46:37 EDT 2011
