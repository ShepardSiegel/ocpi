Bit#(32) compileTime = 1288718619; // Verilog Tue Nov 2 13:23:39 EDT 2010
