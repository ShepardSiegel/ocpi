Bit#(32) compileTime = 1322585792; // Verilog Tue Nov 29 11:56:32 EST 2011
