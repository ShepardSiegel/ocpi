Bit#(32) compileTime = 1289400686; // Verilog Wed Nov 10 09:51:26 EST 2010
