Bit#(32) compileTime = 1295039460; // Verilog Fri Jan 14 16:11:00 EST 2011
