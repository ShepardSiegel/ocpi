<<<<<<< HEAD
Bit#(32) compileTime = 1304787173; // Verilog Sat May 7 12:52:53 EDT 2011
=======
Bit#(32) compileTime = 1304800140; // Verilog Sat May 7 16:29:00 EDT 2011
>>>>>>> 37eff77c6c46b0c0c402ac094217ecdd3d42bd53
