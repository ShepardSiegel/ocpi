Bit#(32) compileTime = 1278684894; // Verilog Fri Jul 9 10:14:54 EDT 2010
