Bit#(32) compileTime = 1279636931; // Verilog Tue Jul 20 10:42:11 EDT 2010
