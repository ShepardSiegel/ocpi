Bit#(32) compileTime = 1328205026; // Verilog Thu Feb 2 12:50:26 EST 2012
