Bit#(32) compileTime = 1276188274; // ISim Thu Jun 10 12:44:34 EDT 2010
