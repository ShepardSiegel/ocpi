Bit#(32) compileTime = 1279898163; // Verilog Fri Jul 23 11:16:03 EDT 2010
