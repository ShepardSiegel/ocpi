Bit#(32) compileTime = 1391543027; // Verilog Tue Feb 4 14:43:47 EST 2014
