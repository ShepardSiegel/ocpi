Bit#(32) compileTime = 1327003947; // Verilog Thu Jan 19 15:12:27 EST 2012
