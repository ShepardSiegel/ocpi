Bit#(32) compileTime = 1275924178; // Verilog Mon Jun 7 11:22:58 EDT 2010
