Bit#(32) compileTime = 1338903437; // Verilog Tue Jun 5 09:37:17 EDT 2012
