Bit#(32) compileTime = 1347452376; // Verilog Wed Sep 12 08:19:36 EDT 2012
