// PCIE.bsv
// Copyright (c) 2009-2012 Atomic Rules LLC - ALL RIGHTS RESERVED

package PCIE;

import PCIEDefs    ::*;  // Types, Functions, and Interfaces
import PCIE_V5     ::*;  // V5 TRN Implementation
import PCIE_V6     ::*;  // V6 TRN Implementation
import PCIE_X6     ::*;  // V6 AXI Implementation
import PCIE_X7     ::*;  // X7 AXI Implementation  (series 7 Xilinx)
import PCIE_S4     ::*;  // S4GX Avalon Implementation

export PCIEDefs    ::*;
export PCIE_V5     ::*;
export PCIE_V6     ::*;
export PCIE_X6     ::*;
export PCIE_X7     ::*;
export PCIE_S4     ::*;

endpackage: PCIE
