Bit#(32) compileTime = 1287149722; // ISim Fri Oct 15 09:35:22 EDT 2010
