Bit#(32) compileTime = 1281619218; // Verilog Thu Aug 12 09:20:18 EDT 2010
