Bit#(32) compileTime = 1292492634; // Verilog Thu Dec 16 04:43:54 EST 2010
