Bit#(32) compileTime = 1279055193; // Verilog Tue Jul 13 17:06:33 EDT 2010
