Bit#(32) compileTime = 1351431278; // Verilog Sun Oct 28 09:34:38 EDT 2012
