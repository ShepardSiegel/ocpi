Bit#(32) compileTime = 1391113942; // Verilog Thu Jan 30 15:32:22 EST 2014
