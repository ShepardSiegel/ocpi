Bit#(32) compileTime = 1299174057; // Verilog Thu Mar 3 12:40:57 EST 2011
