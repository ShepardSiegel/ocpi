Bit#(32) compileTime = 1280524482; // Verilog Fri Jul 30 17:14:42 EDT 2010
