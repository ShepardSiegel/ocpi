Bit#(32) compileTime = 1290111016; // Verilog Thu Nov 18 15:10:16 EST 2010
