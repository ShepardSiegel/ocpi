Bit#(32) compileTime = 1276196525; // Verilog Thu Jun 10 15:02:05 EDT 2010
