Bit#(32) compileTime = 1276702967; // Verilog Wed Jun 16 11:42:47 EDT 2010
