Bit#(32) compileTime = 1287943021; // Verilog Sun Oct 24 13:57:01 EDT 2010
