Bit#(32) compileTime = 1301840560; // Verilog Sun Apr 3 10:22:40 EDT 2011
