Bit#(32) compileTime = 1327784536; // Verilog Sat Jan 28 16:02:16 EST 2012
