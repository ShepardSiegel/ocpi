Bit#(32) compileTime = 1288800604; // Verilog Wed Nov 3 12:10:04 EDT 2010
