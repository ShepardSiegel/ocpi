Bit#(32) compileTime = 1379207501; // Verilog Sat Sep 14 21:11:41 EDT 2013
