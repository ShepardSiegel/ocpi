Bit#(32) compileTime = 1299687790; // Verilog Wed Mar 9 11:23:10 EST 2011
