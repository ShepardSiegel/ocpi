Bit#(32) compileTime = 1281628999; // Verilog Thu Aug 12 12:03:19 EDT 2010
