Bit#(32) compileTime = 1295399918; // Verilog Tue Jan 18 20:18:38 EST 2011
