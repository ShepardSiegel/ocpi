Bit#(32) compileTime = 1290459398; // Verilog Mon Nov 22 15:56:38 EST 2010
