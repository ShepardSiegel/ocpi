Bit#(32) compileTime = 1279113494; // Verilog Wed Jul 14 09:18:14 EDT 2010
