// OCWip.bsv - OpenCPI WIP 
// Copyright (c) 2009-2011 Atomic Rules LLC - ALL RIGHTS RESERVED

package OCWip;

import OCWipDefs    ::*;
import OCPMDefs     ::*;
import OCWci        ::*;
import OCWsi        ::*;
import OCWmi        ::*;
import OCWmemi      ::*;
import OCWti        ::*;

export OCWipDefs    ::*;
export OCPMDefs     ::*;
export OCWci        ::*;
export OCWsi        ::*;
export OCWmi        ::*;
export OCWmemi      ::*;
export OCWti        ::*;


// Cross-Profile Adapter and Convienience IPs...

endpackage: OCWip
