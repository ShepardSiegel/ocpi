Bit#(32) compileTime = 1308584671; // Verilog Mon Jun 20 11:44:31 EDT 2011
