Bit#(32) compileTime = 1292615802; // Verilog Fri Dec 17 14:56:42 EST 2010
