Bit#(32) compileTime = 1289680924; // Verilog Sat Nov 13 15:42:04 EST 2010
