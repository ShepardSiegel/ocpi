Bit#(32) compileTime = 1276264664; // Verilog Fri Jun 11 09:57:44 EDT 2010
