Bit#(32) compileTime = 1278073615; // Verilog Fri Jul 2 08:26:55 EDT 2010
