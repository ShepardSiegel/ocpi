Bit#(32) compileTime = 1328546908; // Verilog Mon Feb 6 11:48:28 EST 2012
