Bit#(32) compileTime = 1284151005; // Verilog Fri Sep 10 16:36:45 EDT 2010
