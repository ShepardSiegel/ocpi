Bit#(32) compileTime = 1286634227; // Verilog Sat Oct 9 10:23:47 EDT 2010
