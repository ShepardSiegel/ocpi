Bit#(32) compileTime = 1304787173; // Verilog Sat May 7 12:52:53 EDT 2011
