Bit#(32) compileTime = 1289910366; // Verilog Tue Nov 16 07:26:06 EST 2010
