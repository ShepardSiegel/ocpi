Bit#(32) compileTime = 1292542626; // Verilog Thu Dec 16 18:37:06 EST 2010
