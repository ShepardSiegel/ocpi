Bit#(32) compileTime = 1288008007; // Bluesim Mon Oct 25 08:00:07 EDT 2010
