Bit#(32) compileTime = 1284377797; // Verilog Mon Sep 13 07:36:37 EDT 2010
