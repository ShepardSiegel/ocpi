// OCWip.bsv - OpenCPI WIP 
// Copyright (c) 2009-2010 Atomic Rules LLC - ALL RIGHTS RESERVED

package OCWip;

import OCWipDefs    ::*;
import OCWci        ::*;
import OCWciOcp     ::*;
import OCWciOcpBfm  ::*;
import OCWciAxi     ::*;
import OCWciAxiBfm  ::*;
import OCWsi        ::*;
import OCWmi        ::*;
import OCWmemi      ::*;
import OCWti        ::*;

export OCWipDefs    ::*;
export OCWci        ::*;
export OCWciOcp     ::*;
export OCWciOcpBfm  ::*;
export OCWciAxi     ::*;
export OCWsi        ::*;
export OCWmi        ::*;
export OCWmemi      ::*;
export OCWti        ::*;


// Cross-Profile Adapter and Convienience IPs...

endpackage: OCWip
