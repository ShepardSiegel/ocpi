Bit#(32) compileTime = 1280260015; // Verilog Tue Jul 27 15:46:55 EDT 2010
