Bit#(32) compileTime = 1290194544; // Verilog Fri Nov 19 14:22:24 EST 2010
