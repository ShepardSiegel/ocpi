Bit#(32) compileTime = 1327972919; // Verilog Mon Jan 30 20:21:59 EST 2012
