Bit#(32) compileTime = 1292500699; // Verilog Thu Dec 16 06:58:19 EST 2010
