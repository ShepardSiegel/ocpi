Bit#(32) compileTime = 1314299939; // Verilog Thu Aug 25 15:18:59 EDT 2011
