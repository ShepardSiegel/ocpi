Bit#(32) compileTime = 1292775325; // Bluesim Sun Dec 19 11:15:25 EST 2010
