Bit#(32) compileTime = 1279021317; // Verilog Tue Jul 13 07:41:57 EDT 2010
