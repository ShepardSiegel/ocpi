Bit#(32) compileTime = 1309030964; // Verilog Sat Jun 25 15:42:44 EDT 2011
