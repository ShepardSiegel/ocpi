Bit#(32) compileTime = 1371848185; // Verilog Fri Jun 21 16:56:25 EDT 2013
