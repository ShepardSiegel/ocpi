Bit#(32) compileTime = 1278417506; // Verilog Tue Jul 6 07:58:26 EDT 2010
