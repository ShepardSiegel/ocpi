Bit#(32) compileTime = 1289737824; // Verilog Sun Nov 14 07:30:24 EST 2010
