Bit#(32) compileTime = 1278772293; // Verilog Sat Jul 10 10:31:33 EDT 2010
