Bit#(32) compileTime = 1297525602; // Verilog Sat Feb 12 10:46:42 EST 2011
