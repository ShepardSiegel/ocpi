Bit#(32) compileTime = 1275847876; // Verilog Sun Jun 6 14:11:16 EDT 2010
