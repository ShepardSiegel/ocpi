Bit#(32) compileTime = 1276792638; // Verilog Thu Jun 17 12:37:18 EDT 2010
