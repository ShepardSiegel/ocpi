Bit#(32) compileTime = 1275662326; // ISim Fri Jun 4 10:38:46 EDT 2010
