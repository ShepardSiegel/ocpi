verilog work ../rtl/lib/BypassWire.v
verilog work ../rtl/lib/SyncFIFO.v
verilog work ../rtl/lib/MakeResetA.v
verilog work ../rtl/lib/SyncResetA.v
verilog work ../rtl/lib/SizedFIFO.v
verilog work ../rtl/lib/FIFO1.v
verilog work ../rtl/lib/FIFO2.v
verilog work ../rtl/lib/RevertReg.v
verilog work ../rtl/lib/BRAM2.v
verilog work ../rtl/lib/BRAM1.v
verilog work ../rtl/lib/BRAM1BE.v
verilog work ../rtl/mkGCDWorker.v
verilog work ../rtl/mkFCAdapter.v
vhdl    work ../vhdl/ocpiTypes.vhd
vhdl    work ../vhdl/biasWorker.vhd
verilog work ../vhdl/mkBiasWorker.v
verilog work ../rtl/mkFPAdapter.v
verilog work ../rtl/mkTLPSM.v
verilog work ../rtl/mkTLPCM.v
verilog work ../rtl/mkPktFork.v
verilog work ../rtl/mkPktMerge.v
verilog work ../rtl/mkOCCP.v
verilog work ../rtl/mkOCDP.v
verilog work ../rtl/mkOCTG.v
verilog work ../rtl/mkOCInf.v
verilog work ../rtl/mkOCApp.v
verilog work ../rtl/mkCTop.v
verilog work ../rtl/mkTB2.v
verilog work ../rtl/lib/main.v

