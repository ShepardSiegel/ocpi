Bit#(32) compileTime = 1276888438; // Verilog Fri Jun 18 15:13:58 EDT 2010
