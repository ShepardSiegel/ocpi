Bit#(32) compileTime = 1286023602; // Verilog Sat Oct 2 08:46:42 EDT 2010
