Bit#(32) compileTime = 1276262115; // Verilog Fri Jun 11 09:15:15 EDT 2010
