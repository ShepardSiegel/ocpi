Bit#(32) compileTime = 1300032374; // Verilog Sun Mar 13 12:06:14 EDT 2011
