Bit#(32) compileTime = 1275410127; // Verilog Tue Jun 1 12:35:27 EDT 2010
