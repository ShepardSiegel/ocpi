<<<<<<< HEAD
Bit#(32) compileTime = 1379207501; // Verilog Sat Sep 14 21:11:41 EDT 2013
=======
Bit#(32) compileTime = 1371848185; // Verilog Fri Jun 21 16:56:25 EDT 2013
>>>>>>> 652a840fab4fae234140a80489c4f89c78f9245c
