Bit#(32) compileTime = 1288362773; // Verilog Fri Oct 29 10:32:53 EDT 2010
