Bit#(32) compileTime = 1295106052; // Verilog Sat Jan 15 10:40:52 EST 2011
