Bit#(32) compileTime = 1294587361; // Verilog Sun Jan 9 10:36:01 EST 2011
