Bit#(32) compileTime = 1355260760; // Verilog Tue Dec 11 16:19:20 EST 2012
