Bit#(32) compileTime = 1289240860; // Verilog Mon Nov 8 13:27:40 EST 2010
