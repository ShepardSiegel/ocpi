Bit#(32) compileTime = 1292688817; // Verilog Sat Dec 18 11:13:37 EST 2010
