Bit#(32) compileTime = 1359067146; // Verilog Thu Jan 24 17:39:06 EST 2013
