Bit#(32) compileTime = 1314185510; // Verilog Wed Aug 24 07:31:50 EDT 2011
