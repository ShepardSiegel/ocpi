Bit#(32) compileTime = 1286722936; // ISim Sun Oct 10 11:02:16 EDT 2010
