Bit#(32) compileTime = 1297287861; // Verilog Wed Feb 9 16:44:21 EST 2011
