Bit#(32) compileTime = 1331051373; // Verilog Tue Mar 6 11:29:33 EST 2012
