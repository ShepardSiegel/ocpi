Bit#(32) compileTime = 1308678764; // Verilog Tue Jun 21 13:52:44 EDT 2011
