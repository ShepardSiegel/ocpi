Bit#(32) compileTime = 1278957614; // Verilog Mon Jul 12 14:00:14 EDT 2010
