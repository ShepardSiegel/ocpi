Bit#(32) compileTime = 1275837022; // Verilog Sun Jun 6 11:10:22 EDT 2010
