Bit#(32) compileTime = 1383230000; // Verilog Thu Oct 31 10:33:20 EDT 2013
