Bit#(32) compileTime = 1359300735; // Verilog Sun Jan 27 10:32:15 EST 2013
