Bit#(32) compileTime = 1289397752; // Verilog Wed Nov 10 09:02:32 EST 2010
