Bit#(32) compileTime = 1288099219; // Bluesim Tue Oct 26 09:20:19 EDT 2010
