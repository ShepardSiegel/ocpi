Bit#(32) compileTime = 1313516659; // Verilog Tue Aug 16 13:44:19 EDT 2011
