Bit#(32) compileTime = 1295106264; // Verilog Sat Jan 15 10:44:24 EST 2011
