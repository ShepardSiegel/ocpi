Bit#(32) compileTime = 1287751220; // Verilog Fri Oct 22 08:40:20 EDT 2010
