Bit#(32) compileTime = 1289393180; // Verilog Wed Nov 10 07:46:20 EST 2010
