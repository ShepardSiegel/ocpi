Bit#(32) compileTime = 1289738647; // Verilog Sun Nov 14 07:44:07 EST 2010
