Bit#(32) compileTime = 1357049537; // Verilog Tue Jan 1 09:12:17 EST 2013
