////////////////////////////////////////////////////////////////////////////////
// Copyright (c) 2009  Bluespec, Inc.   ALL RIGHTS RESERVED.
////////////////////////////////////////////////////////////////////////////////
//  Filename      : Synchronizer.bsv
//  Description   :
////////////////////////////////////////////////////////////////////////////////
package Synchronizer;

// Notes :

////////////////////////////////////////////////////////////////////////////////
/// Imports
////////////////////////////////////////////////////////////////////////////////
import Vector            ::*;

////////////////////////////////////////////////////////////////////////////////
/// Interfaces
////////////////////////////////////////////////////////////////////////////////
(* always_ready, always_enabled *)
interface Synchronizer#(type a);
   method    Action    _write(a x);
   method    a         _read();
endinterface

////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////
///
/// Implementation of Input Synchronizer
///
////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////
module mkSynchronizer#(a initval)(Synchronizer#(a))
   provisos( Bits#(a, sa)
           , Add#(0, sa, 1)
           );

   ////////////////////////////////////////////////////////////////////////////////
   /// Design Elements
   ////////////////////////////////////////////////////////////////////////////////
   Reg#(a)                                   d1                  <- mkReg(initval);
   Reg#(a)                                   d2                  <- mkReg(initval);

   ////////////////////////////////////////////////////////////////////////////////
   /// Interface Connections / Methods
   ////////////////////////////////////////////////////////////////////////////////
   method Action _write(x);
      d1 <= x;
      d2 <= d1;
   endmethod

   method a _read();
      return d2;
   endmethod

endmodule: mkSynchronizer

////////////////////////////////////////////////////////////////////////////////
/// Helper Functions
////////////////////////////////////////////////////////////////////////////////
function Vector#(n,a) readSync(Vector#(n, Synchronizer#(a)) vrin);
   function a readVSync(Synchronizer#(a) i);
      return i._read;
   endfunction
   return map(readVSync, vrin);
endfunction

function Action writeSync(Vector#(n, Synchronizer#(a)) vr, Vector#(n, a) vdin);
   action
      function Action writeVSync(Synchronizer#(a) r, a din);
         action
            r._write(din);
         endaction
      endfunction
      for(Integer i = 0; i < valueof(n); i = i + 1) begin
         writeVSync(vr[i], vdin[i]);
      end
   endaction
endfunction


endpackage: Synchronizer

