Bit#(32) compileTime = 1390768038; // Verilog Sun Jan 26 15:27:18 EST 2014
