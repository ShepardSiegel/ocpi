Bit#(32) compileTime = 1275912093; // Verilog Mon Jun 7 08:01:33 EDT 2010
