// TB10.bsv - A testbench for the PSD
// Copyright (c) 2009-2010 Atomic Rules LLC - ALL RIGHTS RESERVED

import OCWip::*;
import PSD::*;

import Connectable::*;
import GetPut::*;
import Real::*;
import StmtFSM::*;

Bit#(16) tone[64] = {
// Generated by cosgen...
// Freq:64.0000 (samples per radian)
// Freq:0.0312 (fraction of Nyquist)
// Gain:0.9900
  16'h7eb8, // i:   0 phi:0.0000 cosphi:1.0000 
  16'h7e1c, // i:   1 phi:0.0982 cosphi:0.9952 
  16'h7c49, // i:   2 phi:0.1963 cosphi:0.9808 
  16'h7943, // i:   3 phi:0.2945 cosphi:0.9569 
  16'h7513, // i:   4 phi:0.3927 cosphi:0.9239 
  16'h6fc2, // i:   5 phi:0.4909 cosphi:0.8819 
  16'h695d, // i:   6 phi:0.5890 cosphi:0.8315 
  16'h61f5, // i:   7 phi:0.6872 cosphi:0.7730 
  16'h599b, // i:   8 phi:0.7854 cosphi:0.7071 
  16'h5064, // i:   9 phi:0.8836 cosphi:0.6344 
  16'h4667, // i:  10 phi:0.9817 cosphi:0.5556 
  16'h3bbc, // i:  11 phi:1.0799 cosphi:0.4714 
  16'h307e, // i:  12 phi:1.1781 cosphi:0.3827 
  16'h24c9, // i:  13 phi:1.2763 cosphi:0.2903 
  16'h18b9, // i:  14 phi:1.3744 cosphi:0.1951 
  16'h0c6c, // i:  15 phi:1.4726 cosphi:0.0980 
  16'h0000, // i:  16 phi:1.5708 cosphi:-0.0000 
  16'hf395, // i:  17 phi:1.6690 cosphi:-0.0980 
  16'he748, // i:  18 phi:1.7671 cosphi:-0.1951 
  16'hdb38, // i:  19 phi:1.8653 cosphi:-0.2903 
  16'hcf83, // i:  20 phi:1.9635 cosphi:-0.3827 
  16'hc445, // i:  21 phi:2.0617 cosphi:-0.4714 
  16'hb99a, // i:  22 phi:2.1598 cosphi:-0.5556 
  16'haf9d, // i:  23 phi:2.2580 cosphi:-0.6344 
  16'ha666, // i:  24 phi:2.3562 cosphi:-0.7071 
  16'h9e0c, // i:  25 phi:2.4544 cosphi:-0.7730 
  16'h96a4, // i:  26 phi:2.5525 cosphi:-0.8315 
  16'h903f, // i:  27 phi:2.6507 cosphi:-0.8819 
  16'h8aee, // i:  28 phi:2.7489 cosphi:-0.9239 
  16'h86be, // i:  29 phi:2.8471 cosphi:-0.9569 
  16'h83b8, // i:  30 phi:2.9452 cosphi:-0.9808 
  16'h81e5, // i:  31 phi:3.0434 cosphi:-0.9952 
  16'h8149, // i:  32 phi:3.1416 cosphi:-1.0000 
  16'h81e5, // i:  33 phi:3.2398 cosphi:-0.9952 
  16'h83b8, // i:  34 phi:3.3379 cosphi:-0.9808 
  16'h86be, // i:  35 phi:3.4361 cosphi:-0.9569 
  16'h8aee, // i:  36 phi:3.5343 cosphi:-0.9239 
  16'h903f, // i:  37 phi:3.6325 cosphi:-0.8819 
  16'h96a4, // i:  38 phi:3.7306 cosphi:-0.8315 
  16'h9e0c, // i:  39 phi:3.8288 cosphi:-0.7730 
  16'ha666, // i:  40 phi:3.9270 cosphi:-0.7071 
  16'haf9d, // i:  41 phi:4.0252 cosphi:-0.6344 
  16'hb99a, // i:  42 phi:4.1233 cosphi:-0.5556 
  16'hc445, // i:  43 phi:4.2215 cosphi:-0.4714 
  16'hcf83, // i:  44 phi:4.3197 cosphi:-0.3827 
  16'hdb38, // i:  45 phi:4.4179 cosphi:-0.2903 
  16'he748, // i:  46 phi:4.5160 cosphi:-0.1951 
  16'hf395, // i:  47 phi:4.6142 cosphi:-0.0980 
  16'h0000, // i:  48 phi:4.7124 cosphi:0.0000 
  16'h0c6c, // i:  49 phi:4.8106 cosphi:0.0980 
  16'h18b9, // i:  50 phi:4.9087 cosphi:0.1951 
  16'h24c9, // i:  51 phi:5.0069 cosphi:0.2903 
  16'h307e, // i:  52 phi:5.1051 cosphi:0.3827 
  16'h3bbc, // i:  53 phi:5.2033 cosphi:0.4714 
  16'h4667, // i:  54 phi:5.3014 cosphi:0.5556 
  16'h5064, // i:  55 phi:5.3996 cosphi:0.6344 
  16'h599b, // i:  56 phi:5.4978 cosphi:0.7071 
  16'h61f5, // i:  57 phi:5.5960 cosphi:0.7730 
  16'h695d, // i:  58 phi:5.6941 cosphi:0.8315 
  16'h6fc2, // i:  59 phi:5.7923 cosphi:0.8819 
  16'h7513, // i:  60 phi:5.8905 cosphi:0.9239 
  16'h7943, // i:  61 phi:5.9887 cosphi:0.9569 
  16'h7c49, // i:  62 phi:6.0868 cosphi:0.9808 
  16'h7e1c  // i:  63 phi:6.1850 cosphi:0.9952 
};

(* synthesize *)
module mkTB10();

  Reg#(Bit#(16))              simCycle       <- mkReg(0);       // simulation cycle counter
  WciEMasterIfc#(20,32)       wci            <- mkWciEMaster;    // WCI-OCP-Master convienenice logic
  WsiMasterIfc#(12,32,4,8,0)  wsiM           <- mkWsiMaster;    // WSI-OCP-Master convienenice logic
  WsiSlaveIfc #(12,32,4,8,0)  wsiS           <- mkWsiSlave;     // WSI-OCP-Slave  convienenice logic

  // It is each WCI master's job to generate for each WCI M-S pairing a mReset_n signal that can reset each worker
  // We send that reset in on the "reset_by" line to reset all state associated with worker module...
  PSDIfc                      psdWorker      <- mkPSD(32'h00000000, True, reset_by wci.mas.mReset_n);   // instance the PSD DUT

  Reg#(Bool)                  enWsiSource    <- mkReg(False);   // Trigger for WSI generator
  Reg#(Bool)                  enWsiChecker   <- mkReg(False);   // Trigger for WSI checker
  Reg#(Bool)                  testOperating  <- mkReg(False);   // Enable for test Operating
  Reg#(Bit#(16))              srcMesgCount   <- mkReg(0);       // Number of Messages sent
  Reg#(Bit#(16))              srcUnrollCnt   <- mkReg(0);       // Message Positions to go
  Reg#(Bit#(32))              srcDataOut     <- mkReg(0);       // DWORD ordinal count
  Reg#(Bit#(6))               srcIndex       <- mkReg(0);       // Src Tone Index
  Reg#(Bit#(16))              dstMesgCount   <- mkReg(0);       // Number of Messages sent
  Reg#(Bit#(16))              dstUnrollCnt   <- mkReg(0);       // Message Positions to go
  Reg#(Bit#(32))              dstDataOut     <- mkReg(0);       // DWORD ordinal count

  mkConnection(wci.mas,  psdWorker.wciS0);             // connect the WCI Master to the DUT
  mkConnection(toWsiEM(wsiM.mas), psdWorker.wsiS0);    // connect the Source wsiM to the psdWorker wsi-S input
  Wsi_Es#(12,32,4,8,0) wsi_Es <- mkWsiStoES(wsiS.slv); // Convert the conventional to explicit 
  mkConnection(psdWorker.wsiM0,  wsi_Es);              // connect the psdWorker wsi-M output to the Sinc wsiS

  // WCI Interaction
  // A sequence of control-configuration operartions to be performed...
  Stmt wciSeq = 
  seq
    $display("[%0d]: %m: Checking for DUT presence...", $time);
    await(wci.present);

    $display("[%0d]: %m: Taking DUT out of Reset...", $time);
    wci.req(Admin, True,  20'h00_0024, 'h8000_0004, 'hF);
    action let r <- wci.resp; endaction

    $display("[%0d]: %m: CONTROL-OP: -INITIALIZE- DUT...", $time);
    wci.req(Control, False, 20'h00_0000, ?, ?);
    action let r <- wci.resp; endaction

    $display("[%0d]: %m: Write Dataplane Config Properties...", $time);
    wci.req(Config, True, 20'h00_0004, 32'h0000_0002, 'hF);                     // psdCtrl
    action let r <- wci.resp; endaction

    $display("[%0d]: %m: Read Dataplane Config Properties...", $time);
    wci.req(Config, False, 20'h00_0004, ?, ?);
    action let r <- wci.resp; endaction

    $display("[%0d]: %m: CONTROL-OP: -START- DUT...", $time);
    wci.req(Control, False, 20'h00_0004, ?, ?);
    action let r <- wci.resp; endaction

    testOperating <= True;
    dstUnrollCnt  <= 2048;
    enWsiChecker  <= True;

    srcUnrollCnt  <= 2048;
    enWsiSource   <= True;
  endseq;
  FSM  wciSeqFsm  <- mkFSM(wciSeq);
  Once wciSeqOnce <- mkOnce(wciSeqFsm.start);

  // Start of the WCI sequence...
  rule runWciSeq;
    wciSeqOnce.start;
  endrule

  // This rule inhibits dataflow on the WSI ports until the WCI port isOperating...
  rule operating_actions (testOperating);
    wsiS.operate();
    wsiM.operate();
  endrule

  // WSI Interaction
  // Producer Stream...
  rule wsi_source (enWsiSource);
    Bool lastWord  = (srcUnrollCnt == 1);
    Bit#(8) opcode = 0;
    Bit#(16) wsiBurstLength = 2048; // in Words (4B)

    if (srcMesgCount < 1)
      wsiM.reqPut.put (WsiReq    {cmd  : WR ,
                               reqLast : lastWord,
                               reqInfo : opcode,
                          burstPrecise : False,
                           burstLength : '1,
                               //data  : {srcDataOut[15:0],srcDataOut[15:0]},
                                 data  : {tone[srcIndex+1],tone[srcIndex]},
                               byteEn  : '1,
                             dataInfo  : '0 });

    srcIndex <= srcIndex + 2;
    srcDataOut  <= srcDataOut  + 1;
    if (lastWord) begin
      srcMesgCount <= srcMesgCount + 1;
      $display("[%0d]: %m: wsi_source: End of WSI Producer Egress: srcMesgCount:%0x opcode:%0x", $time, srcMesgCount, opcode);
    end
    srcUnrollCnt <= (lastWord) ? wsiBurstLength : srcUnrollCnt - 1;
  endrule

  // Consume Stream...
  rule wsi_checker (enWsiChecker);
    Bit#(8) opcode = wsiS.reqPeek.reqInfo;
    Bit#(16) wsiBurstLength =  extend(wsiS.reqPeek.burstLength);
    Bit#(16) mesgLengthB    =  wsiBurstLength<<2;
    Bool lastWord  = (dstUnrollCnt == 1);
    WsiReq#(12,32,4,8,0) w <- wsiS.reqGet.get;

    Bit#(32) dataGot = w.data;

    //Bit#(32) dataExp = dstDataOut;
    //if (dataGot != dataExp) $display("[%0d]: %m: wsi_checker MISMATCH: exp:%0x got:%0x srcMesgCount:%0x", $time, dataExp, dataGot, dstMesgCount);

    $display("[%0d]: %m: PSD bin:%0d %04x, bin:%0d %04x", $time, dstDataOut, dataGot[15:0], dstDataOut+1, dataGot[31:16]);

    dstDataOut  <= dstDataOut  + 2;
    if (lastWord) begin
      dstMesgCount <= dstMesgCount + 1;
      $display("[%0d]: %m: wsi_source: End of WSI Consumer Ingress: dstMesgCount:%0x opcode:%0x", $time, dstMesgCount, opcode);
    end
    dstUnrollCnt <= (lastWord) ? wsiBurstLength : dstUnrollCnt - 1;
  endrule

  // Simulation Control...
  rule increment_simCycle;
    simCycle <= simCycle + 1;
  endrule

  rule terminate (simCycle==20000);
    $display("[%0d]: %m: mkTB10 termination", $time);
    $finish;
  endrule

endmodule: mkTB10

