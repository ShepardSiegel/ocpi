Bit#(32) compileTime = 1281639883; // Verilog Thu Aug 12 15:04:43 EDT 2010
