Bit#(32) compileTime = 1304954458; // Verilog Mon May 9 11:20:58 EDT 2011
