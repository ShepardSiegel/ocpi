Bit#(32) compileTime = 1281526382; // Verilog Wed Aug 11 07:33:02 EDT 2010
