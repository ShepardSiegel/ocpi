Bit#(32) compileTime = 1295466944; // Verilog Wed Jan 19 14:55:44 EST 2011
