Bit#(32) compileTime = 1354117072; // Verilog Wed Nov 28 10:37:52 EST 2012
