Bit#(32) compileTime = 1279897561; // Verilog Fri Jul 23 11:06:01 EDT 2010
