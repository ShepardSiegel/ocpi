Bit#(32) compileTime = 1302556156; // Verilog Mon Apr 11 17:09:16 EDT 2011
