Bit#(32) compileTime = 1296079549; // Verilog Wed Jan 26 17:05:49 EST 2011
