Bit#(32) compileTime = 1288043992; // Verilog Mon Oct 25 17:59:52 EDT 2010
