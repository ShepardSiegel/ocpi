Bit#(32) compileTime = 1278786937; // Verilog Sat Jul 10 14:35:37 EDT 2010
