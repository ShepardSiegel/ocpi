Bit#(32) compileTime = 1296837410; // Verilog Fri Feb 4 11:36:50 EST 2011
