Bit#(32) compileTime = 1277295491; // Verilog Wed Jun 23 08:18:11 EDT 2010
