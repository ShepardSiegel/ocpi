Bit#(32) compileTime = 1379248177; // Verilog Sun Sep 15 08:29:37 EDT 2013
