Bit#(32) compileTime = 1288735921; // Verilog Tue Nov 2 18:12:01 EDT 2010
