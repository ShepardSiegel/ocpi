Bit#(32) compileTime = 1278844952; // Verilog Sun Jul 11 06:42:32 EDT 2010
