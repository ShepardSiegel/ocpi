Bit#(32) compileTime = 1281462596; // Verilog Tue Aug 10 13:49:56 EDT 2010
