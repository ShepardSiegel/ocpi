Bit#(32) compileTime = 1292527182; // Verilog Thu Dec 16 14:19:42 EST 2010
