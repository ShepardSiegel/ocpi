Bit#(32) compileTime = 1330533871; // Verilog Wed Feb 29 11:44:31 EST 2012
