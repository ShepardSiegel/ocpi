Bit#(32) compileTime = 1297282035; // Bluesim Wed Feb 9 15:07:15 EST 2011
