Bit#(32) compileTime = 1351436476; // Verilog Sun Oct 28 11:01:16 EDT 2012
