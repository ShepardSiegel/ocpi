Bit#(32) compileTime = 1383162921; // Verilog Wed Oct 30 15:55:21 EDT 2013
