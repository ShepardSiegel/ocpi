Bit#(32) compileTime = 1282230022; // Verilog Thu Aug 19 11:00:22 EDT 2010
