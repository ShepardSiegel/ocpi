Bit#(32) compileTime = 1303937181; // Verilog Wed Apr 27 16:46:21 EDT 2011
