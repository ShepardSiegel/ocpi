Bit#(32) compileTime = 1330523962; // Verilog Wed Feb 29 08:59:22 EST 2012
