Bit#(32) compileTime = 1278945858; // Verilog Mon Jul 12 10:44:18 EDT 2010
