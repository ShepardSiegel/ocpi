Bit#(32) compileTime = 1276177455; // ISim Thu Jun 10 09:44:15 EDT 2010
