Bit#(32) compileTime = 1325689641; // Verilog Wed Jan 4 10:07:21 EST 2012
