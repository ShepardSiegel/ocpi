Bit#(32) compileTime = 1331046544; // Verilog Tue Mar 6 10:09:04 EST 2012
