// ARAXI.bsv - The Atomic Rules AXI Packages 
// Copyright (c) 2009-2011 Atomic Rules LLC - ALL RIGHTS RESERVED

package ARAXI;

import ARAXI4L    ::*;  // AXI4-Lite   (A4L)
import ARAXI4S    ::*;  // AXI4-Stream (AXIS)

export ARAXI4L    ::*;
export ARAXI4S    ::*;

endpackage: ARAXI
