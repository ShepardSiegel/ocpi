Bit#(32) compileTime = 1276800010; // Verilog Thu Jun 17 14:40:10 EDT 2010
