Bit#(32) compileTime = 1383146627; // Verilog Wed Oct 30 11:23:47 EDT 2013
