Bit#(32) compileTime = 1277139201; // Verilog Mon Jun 21 12:53:21 EDT 2010
