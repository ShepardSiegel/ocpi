Bit#(32) compileTime = 1308858805; // Verilog Thu Jun 23 15:53:25 EDT 2011
