Bit#(32) compileTime = 1391459380; // Verilog Mon Feb 3 15:29:40 EST 2014
