Bit#(32) compileTime = 1280189777; // Verilog Mon Jul 26 20:16:17 EDT 2010
