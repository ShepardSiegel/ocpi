Bit#(32) compileTime = 1281628055; // Verilog Thu Aug 12 11:47:35 EDT 2010
