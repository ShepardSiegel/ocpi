Bit#(32) compileTime = 1314645303; // Verilog Mon Aug 29 15:15:03 EDT 2011
