Bit#(32) compileTime = 1306183624; // Verilog Mon May 23 16:47:04 EDT 2011
