Bit#(32) compileTime = 1288807307; // Verilog Wed Nov 3 14:01:47 EDT 2010
