Bit#(32) compileTime = 1289218332; // Verilog Mon Nov 8 07:12:12 EST 2010
