Bit#(32) compileTime = 1287065510; // Verilog Thu Oct 14 10:11:50 EDT 2010
