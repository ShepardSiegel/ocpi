Bit#(32) compileTime = 1277481406; // Verilog Fri Jun 25 11:56:46 EDT 2010
