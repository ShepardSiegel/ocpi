Bit#(32) compileTime = 1275943709; // Verilog Mon Jun 7 16:48:29 EDT 2010
