Bit#(32) compileTime = 1275426555; // Verilog Tue Jun 1 17:09:15 EDT 2010
