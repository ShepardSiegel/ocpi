Bit#(32) compileTime = 1281704041; // Verilog Fri Aug 13 08:54:01 EDT 2010
