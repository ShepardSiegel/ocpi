Bit#(32) compileTime = 1337778735; // Verilog Wed May 23 09:12:15 EDT 2012
