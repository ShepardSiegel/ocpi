Bit#(32) compileTime = 1289252933; // Verilog Mon Nov 8 16:48:53 EST 2010
