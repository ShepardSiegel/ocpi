Bit#(32) compileTime = 1286322778; // Verilog Tue Oct 5 19:52:58 EDT 2010
