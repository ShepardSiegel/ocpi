Bit#(32) compileTime = 1277999220; // Verilog Thu Jul 1 11:47:00 EDT 2010
