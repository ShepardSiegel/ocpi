Bit#(32) compileTime = 1281708527; // Verilog Fri Aug 13 10:08:47 EDT 2010
