Bit#(32) compileTime = 1321968593; // Verilog Tue Nov 22 08:29:53 EST 2011
