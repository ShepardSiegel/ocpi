Bit#(32) compileTime = 1283192366; // ISim Mon Aug 30 14:19:26 EDT 2010
