Bit#(32) compileTime = 1383673480; // Verilog Tue Nov 5 12:44:40 EST 2013
