// UUID generated for platform 'n210', device '(null)', uuid '2aa339ca-c822-4067-9c4c-d943f3195a48'
module mkUUID(uuid);
output [511 : 0] uuid;
wire [511 : 0] uuid = 512'haeaee44f2aa339cac82240679c4cd943f3195a486e3231300000000000000000000000007863337364333430306100000000000000000000b9d7400000000000;
endmodule // mkUUID
