Bit#(32) compileTime = 1288469489; // Verilog Sat Oct 30 16:11:29 EDT 2010
