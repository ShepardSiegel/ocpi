Bit#(32) compileTime = 1276036878; // Verilog Tue Jun 8 18:41:18 EDT 2010
