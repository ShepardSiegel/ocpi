Bit#(32) compileTime = 1304800140; // Verilog Sat May 7 16:29:00 EDT 2011
