Bit#(32) compileTime = 1276710388; // Verilog Wed Jun 16 13:46:28 EDT 2010
