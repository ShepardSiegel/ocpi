Bit#(32) compileTime = 1327005233; // Verilog Thu Jan 19 15:33:53 EST 2012
