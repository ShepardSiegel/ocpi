Bit#(32) compileTime = 1390838362; // Verilog Mon Jan 27 10:59:22 EST 2014
