Bit#(32) compileTime = 1323201679; // Verilog Tue Dec 6 15:01:19 EST 2011
