Bit#(32) compileTime = 1292511991; // Verilog Thu Dec 16 10:06:31 EST 2010
