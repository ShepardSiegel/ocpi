Bit#(32) compileTime = 1279649143; // Verilog Tue Jul 20 14:05:43 EDT 2010
