Bit#(32) compileTime = 1304782851; // Verilog Sat May 7 11:40:51 EDT 2011
