Bit#(32) compileTime = 1279997335; // Verilog Sat Jul 24 14:48:55 EDT 2010
